module BCD_to_7seg (
    input [4:0] BCD,
    output [6:0] seg
);
    always @(*) begin
        case(BCD)
            5'b00000: seg = 7'b0111111; // 0
            5'b00001: seg = 7'b0000110; // 1
            5'b00010: seg = 7'b1011011; // 2
            5'b00011: seg = 7'b1001111; // 3
            5'b00100: seg = 7'b1100110; // 4
            5'b00101: seg = 7'b1101101; // 5
            5'b00110: seg = 7'b1111101; // 6
            5'b00111: seg = 7'b0000111; // 7
            5'b01000: seg = 7'b1111111; // 8
            5'b01001: seg = 7'b1101111; // 9
            5'b01010: seg = 7'b1110111; // 10
            5'b01011: seg = 7'b1111110; // 11
            5'b01100: seg = 7'b0111001; // 12
            5'b01101: seg = 7'b1011111; // 13
            5'b01110: seg = 7'b1111001; // 14
            5'b01111: seg = 7'b1110000; // 15
            5'b10000: seg = 7'b1111111; // 16
            5'b10001: seg = 7'b0000110; // 17
            5'b10010: seg = 7'b1011011; // 18
            5'b10011: seg = 7'b1001111; // 19
            default:  seg = 7'b0000000; 
        endcase
    end
endmodule
